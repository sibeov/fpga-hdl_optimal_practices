-- Standard IEEE library.
library ieee;
context ieee.ieee_std_context;

entity bare_entity is
	generic (
		-- Generics
	);
	port (
		-- Physical ports
	);
end entity bare_entity;

architecture rtl of bare_entity is

	-- Declarative section of architecture

begin

	-- Concurrent section of architecture

end architecture rtl;